`timescale 1ns / 1ps



//Percent Effort
// Roes: 33% Evan: 33% Noah: 33%
////////////////////////////////////////////////////////////////////////////////
// ECE369A - Computer Architecture
// Laboratory  
// Module - PCAdder.v
// Description - 32-Bit program counter (PC) adder.
// 
// INPUTS:-
// PCResult: 32-Bit input port.
// 
// OUTPUTS:-
// PCAddResult: 32-Bit output port.
//
// FUNCTIONALITY:-
// Design an incrementor (or a hard-wired ADD ALU whose first input is from the 
// PC, and whose second input is a hard-wired 4) that computes the current 
// PC + 4. The result should always be an increment of the signal 'PCResult' by 
// 4 (i.e., PCAddResult = PCResult + 4).
////////////////////////////////////////////////////////////////////////////////

module PCAdder(PCResult, PCAddResult);

    input [31:0] PCResult;          // Current PC value coming from ProgramCounter
    output[31:0] PCAddResult;  // Next PC value (PC + 4), fed back into ProgramCounter

    assign PCAddResult = PCResult + 4; // Increment the PC by 4 (word-aligned instruction step)
  
    /* The logic is complete here:
       - This is essentially a hard-wired adder.
       - Every instruction in MIPS is 4 bytes, so we increment PC by 4 each time.
       - PCAddResult is then fed back to ProgramCounter in the Instruction Fetch Unit. */
endmodule

