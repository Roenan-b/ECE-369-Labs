`timescale 1ns / 1ps

module AND(A, B, out);

  input A;
  input B;
  output out;

  assign out = A & B;

endmodule
