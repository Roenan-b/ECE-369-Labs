`timescale 1ns / 1ps


module RegisterID_EX(ReadData1In, ReadData1Out, ReadData2In, ReadData2Out,
                     Instruction1In, Instruction1Out, Instruction2In, Instruction2Out, Instruction3In, Instruction3Out, 
