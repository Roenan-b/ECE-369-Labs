module immSL2(in, out);
